interface add_if;
  logic clk;
  logic reset;
  logic [7:0] in1;
  logic [7:0] in2;
  logic [8:0] out;
  
endinterface
